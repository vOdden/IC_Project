[aimspice]
[description]
1842
* Simulation of one pixel


.include C:\Users\sigur\OneDrive\Skrivebord\DIC_Project\p18_cmos_models_tt.inc
!.include p18_model_card.inc

*
*	Parameters
*
.param L1 = 1.08u
.param W1 = 1.08u
.param L2 = 1.08u
.param W2 = 1.08u
.param L3 = 0.67u
.param W3 = 3.00u
.param L4 = 1.08u
.param W4 = 5.04u
.param MCL = 0.36u
.param MCW = 5.04u
.param CSvalue = 2pF
.param CCvalue = 3pF
*
*	Circuitry
*
XPD1 Vdd N1 PhotoDiode
MN1 N1 Expose N2 0 NMOS L=L1 W=W1
MN2 N2 Erase 0 0 NMOS L=L2 W=W2
CS N2 0 CSvalue
MP3 0 N2 N3 Vdd PMOS L=L3 W=W3
MP4 N3 NRE Out Vdd PMOS L=L4 W=W4

MC Out Out Vdd Vdd PMOS L=MCL W=MCW
CC Out 0 CCvalue

*
*	Testbench
*
.param Ipd_1 = 750p ! Photodiode current, [50pA, 750pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 2m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

VDD Vdd 0 dc VDD
VEXPOSE Expose 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE Erase 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE NRE 0 dc 0 pulse(VDD 0 NRE_DLY TRF TRF CLK_PERIOD PERIOD)

.plot V(EXPOSE) V(ERASE) V(NRE) V(Out) V(N2) V(N3)
.plot V(out)

*
*	PHOTODIODE 
*
.subckt PhotoDiode  VDD N1_R1C1
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1
d1 N1_R1C1 vdd dwell 1
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40
Cd1 N1_R1C1 VDD 30f
.ends 
[dc]
1
I1_R1C1
0
5
0.01
[tran]
0.1
60ms
X
X
0
[ana]
4 1
0
1 1
1 1 -0.5 2
3
v(n1)
v(n2)
v(n3)
[end]
