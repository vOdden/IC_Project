[aimspice]
[description]
1889
*	One pixel


.include C:\Users\sigur\OneDrive\Skrivebord\DIC_Project\p18_cmos_models_tt.inc
!.include C:\Users\sigur\OneDrive\Skrivebord\DIC_v2\p18_model_card.inc

.param Ipd_1 = 750p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 2m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal


VDD Vdd 0 dc VDD
*X1 Vdd 0 EXPOSE ERASE Out Exposecircuit
X2 Vdd 0 Expose Erase NRE Out OnePixel


VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE NRE 0 dc 0 pulse(VDD 0 NRE_DLY TRF TRF CLK_PERIOD PERIOD)

.plot V(EXPOSE) V(ERASE) V(NRE) V(Out)
*.plot V(Out)


.subckt OnePixel Vdd Vss Expose Erase NRE Out
XExp Vdd Vss Expose Erase N2 Exposecircuit
MP3 Vss N2 N3 Vdd PMOS L=1u W=5u
MP4 N3 NRE Out Vdd PMOS L=0.7u W=10u
*Xload Vdd Vss Out LoadTransistor

.ends

.subckt LoadTransistor Vdd Vss Gate
MC Gate Gate Vdd Vdd PMOS L=2u W=10u
CC Gate Vss 3p
.ends

.subckt Exposecircuit Vdd Vss Expose Erase N2
XPD1 Vdd N1 PhotoDiode
MN1 N1 Expose N2 Vss NMOS L=0.7u W=10u
MN2 N2 Erase Vss Vss NMOS L=2u W=2u
CS N2 Vss 1.5p
.ends

.subckt PhotoDiode  VDD N1_R1C1
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1
d1 N1_R1C1 vdd dwell 1
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40
Cd1 N1_R1C1 VDD 30f
.ends 
[dc]
1
VDD
0
1
0.001
[ana]
1 0
[end]
