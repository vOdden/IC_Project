[aimspice]
[description]
2288
*	All four pixels

.include C:\Users\sigur\OneDrive\Skrivebord\DIC_Project\p18_cmos_models_tt.inc

*
*	Parameters
*
.param L1 = 0.7u
.param W1 = 3u
.param L2 = 0.7u
.param W2 = 3u
.param L3 = 1.08u
.param W3 = 5.04u
.param L4 = 1.08u		!
.param W4 = 5.04u		!
.param MCL = 1.08u 	!
.param MCW = 5.04u	!
.param CSvalue = 1.5pF	!
.param CCvalue = 3pF	!

XONEPIXEL11 VDD 0 Expose Erase NRE_R1 OUT1 OnePixel
XONEPIXEL12 VDD 0 Expose Erase NRE_R1 OUT2 OnePixel
XONEPIXEL21 VDD 0 Expose Erase NRE_R2 OUT1 OnePixel
XONEPIXEL22 VDD 0 Expose Erase NRE_R2 OUT2 OnePixel

*
*	Testbench
*
.param Ipd_1 = 50p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 30m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE signal
.param NRE_R2_DLY = {4*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

VDD Vdd 0 dc VDD
VEXPOSE Expose 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE Erase 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R1 NRE_R1 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R2 NRE_R2 0 dc 0 pulse(VDD 0 NRE_R2_DLY TRF TRF CLK_PERIOD PERIOD)

.plot V(EXPOSE) V(ERASE) V(Out1) V(Out2) V(NRE_R1) V(NRE_R2)
.plot V(Out1) V(Out2)
.plot V(NRE_R1) V(NRE_R2) V(N2)

*
*	One Pixel circuit
*

.subckt OnePixel Vdd Vss Expose Erase NRE Out
XPD1 Vdd N1 PhotoDiode
MN1 N1 Expose N2 0 NMOS L=L1 W=W1
MN2 N2 Erase 0 0 NMOS L=L2 W=W2
CS N2 0 CSvalue
MP3 0 N2 N3 Vdd PMOS L=L3 W=W3
MP4 N3 NRE Out Vdd PMOS L=L4 W=W4

MC Out Out Vdd Vdd PMOS L=MCL W=MCW
CC Out 0 CCvalue
.ends

.subckt PhotoDiode  VDD N1_R1C1
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1
d1 N1_R1C1 vdd dwell 1
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40
Cd1 N1_R1C1 VDD 30f
.ends
[dc]
1
I1_R1C1
0
5
0.01
[tran]
0.01
60ms
X
X
0
[ana]
4 0
[end]
